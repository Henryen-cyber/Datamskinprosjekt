`include "types.sv"

module RayTraceDatapath (
    input logic       clk,
    input logic[1:0]  index,
    output logic      valid
    );

    always @(posedge clk) begin
        
    end    

endmodule
