`include "in_spi.sv"
`include "bind_spi.sv"
module tb();

    in_spi uin_spi();

endmodule
