program testPr_spi(
    in_spi uin_spi
);

//Implement tasks and immediate assertions

endprogram

